module mux_tb;

endmodule;